// command line for phase debug: +access+r +UVM_PHASE_TRACE
// command line for objection debug: +access+r +UVM_OBJECTION_TRACE
